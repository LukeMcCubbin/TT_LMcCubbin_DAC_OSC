magic
tech sky130A
timestamp 1698067942
<< pwell >>
rect -557 -369 557 369
<< psubdiff >>
rect -539 334 539 351
rect -539 -334 -522 334
rect 522 -334 539 334
rect -539 -351 -491 -334
rect 491 -351 539 -334
<< psubdiffcont >>
rect -491 -351 491 -334
<< xpolycontact >>
rect -474 70 -439 286
rect -474 -286 -439 -70
rect -391 70 -356 286
rect -391 -286 -356 -70
rect -308 70 -273 286
rect -308 -286 -273 -70
rect -225 70 -190 286
rect -225 -286 -190 -70
rect -142 70 -107 286
rect -142 -286 -107 -70
rect -59 70 -24 286
rect -59 -286 -24 -70
rect 24 70 59 286
rect 24 -286 59 -70
rect 107 70 142 286
rect 107 -286 142 -70
rect 190 70 225 286
rect 190 -286 225 -70
rect 273 70 308 286
rect 273 -286 308 -70
rect 356 70 391 286
rect 356 -286 391 -70
rect 439 70 474 286
rect 439 -286 474 -70
<< xpolyres >>
rect -474 -70 -439 70
rect -391 -70 -356 70
rect -308 -70 -273 70
rect -225 -70 -190 70
rect -142 -70 -107 70
rect -59 -70 -24 70
rect 24 -70 59 70
rect 107 -70 142 70
rect 190 -70 225 70
rect 273 -70 308 70
rect 356 -70 391 70
rect 439 -70 474 70
<< locali >>
rect -499 -351 -491 -334
rect 491 -351 499 -334
<< properties >>
string FIXED_BBOX -530 -342 530 342
<< end >>
