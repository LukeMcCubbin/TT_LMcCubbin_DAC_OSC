magic
tech sky130A
magscale 1 2
timestamp 1760635213
use sky130_fd_pr__res_xhigh_po_0p35_KD7KM5  sky130_fd_pr__res_xhigh_po_0p35_KD7KM5_0
timestamp 1760635213
transform 1 0 729 0 1 579
box -782 -632 782 632
<< end >>
