magic
tech sky130A
magscale 1 2
timestamp 1759518956
<< error_p >>
rect 4227 -1371 4280 -1370
rect 4209 -1405 4280 -1371
rect 4210 -1406 4280 -1405
rect 4227 -1440 4298 -1406
rect 1131 -3181 1166 -3164
rect 1132 -3182 1166 -3181
rect 1132 -3218 1202 -3182
rect 1149 -3252 1220 -3218
rect 1149 -3613 1219 -3252
rect 1149 -3649 1202 -3613
rect 3490 -3666 3505 -3218
rect 3524 -3666 3558 -3164
rect 3524 -3700 3539 -3666
rect 4227 -3719 4297 -1440
rect 4949 -3341 4983 -3323
rect 7341 -3341 7375 -3323
rect 4949 -3377 5019 -3341
rect 4966 -3411 5037 -3377
rect 4227 -3755 4280 -3719
rect 4966 -3772 5036 -3411
rect 4966 -3808 5019 -3772
rect 7305 -3825 7375 -3341
rect 7305 -3861 7358 -3825
rect 4107 -7959 4160 -7958
rect 4089 -7993 4160 -7959
rect 4090 -7994 4160 -7993
rect 4107 -8028 4178 -7994
rect 1011 -9769 1046 -9752
rect 1012 -9770 1046 -9769
rect 1012 -9806 1082 -9770
rect 1029 -9840 1100 -9806
rect 1029 -10201 1099 -9840
rect 1029 -10237 1082 -10201
rect 3370 -10254 3385 -9806
rect 3404 -10254 3438 -9752
rect 3404 -10288 3419 -10254
rect 4107 -10307 4177 -8028
rect 4829 -9929 4863 -9911
rect 7221 -9929 7255 -9911
rect 4829 -9965 4899 -9929
rect 4846 -9999 4917 -9965
rect 4107 -10343 4160 -10307
rect 4846 -10360 4916 -9999
rect 4846 -10396 4899 -10360
rect 7185 -10413 7255 -9929
rect 7185 -10449 7238 -10413
rect 3957 -14409 4010 -14408
rect 3939 -14443 4010 -14409
rect 3940 -14444 4010 -14443
rect 3957 -14478 4028 -14444
rect 861 -16219 896 -16202
rect 862 -16220 896 -16219
rect 862 -16256 932 -16220
rect 879 -16290 950 -16256
rect 879 -16651 949 -16290
rect 879 -16687 932 -16651
rect 3220 -16704 3235 -16256
rect 3254 -16704 3288 -16202
rect 3254 -16738 3269 -16704
rect 3957 -16757 4027 -14478
rect 4679 -16379 4713 -16361
rect 7071 -16379 7105 -16361
rect 4679 -16415 4749 -16379
rect 4696 -16449 4767 -16415
rect 3957 -16793 4010 -16757
rect 4696 -16810 4766 -16449
rect 4696 -16846 4749 -16810
rect 7035 -16863 7105 -16379
rect 7035 -16899 7088 -16863
<< metal1 >>
rect -6062 -362 -5862 -162
rect -6062 -762 -5862 -562
rect -6062 -1162 -5862 -962
rect -6062 -1562 -5862 -1362
use ringosc_buf  xbuf1
timestamp 1759517325
transform 1 0 -6900 0 1 -3986
box 1170 -506 4008 2030
use ringosc_buf  xbuf2
timestamp 1759517325
transform 1 0 -6976 0 1 -14764
box 1170 -506 4008 2030
use ringosc_buf  xbuf3
timestamp 1759517325
transform 1 0 -6938 0 1 -9450
box 1170 -506 4008 2030
use ringosc_delay  xro1
timestamp 1759517188
transform 1 0 -1098 0 1 -7630
box -212 -2872 8875 2090
use ringosc_delay  xro2
timestamp 1759517188
transform 1 0 -1248 0 1 -14080
box -212 -2872 8875 2090
use ringosc_delay  xro3
timestamp 1759517188
transform 1 0 -978 0 1 -1042
box -212 -2872 8875 2090
<< labels >>
flabel metal1 -6062 -1562 -5862 -1362 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 -6062 -1162 -5862 -962 0 FreeSans 256 0 0 0 ena
port 2 nsew
flabel metal1 -6062 -762 -5862 -562 0 FreeSans 256 0 0 0 clk_out
port 1 nsew
flabel metal1 -6062 -362 -5862 -162 0 FreeSans 256 0 0 0 vdd
port 0 nsew
<< end >>
