** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/tt_um_tt05_analog_test_combined.sch
.subckt tt_um_tt05_analog_test_combined uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] VPWR
+ uio_out[0] uio_out[1] clk uio_out[2] ena rst_n uio_out[3] uio_out[4] uio_out[5] uio_out[6] ui_in[0] ui_in[1] uio_out[7] ui_in[2] uo_out[0]
+ ui_in[3] uo_out[1] ui_in[4] ui_in[5] uo_out[2] ui_in[6] uo_out[3] ui_in[7] uo_out[4] uo_out[5] uio_in[0] uo_out[6] uio_in[1] uo_out[7]
+ uio_in[2] uio_in[3] ua[0] uio_in[4] ua[1] uio_in[5] ua[2] uio_in[6] ua[3] uio_in[7] ua[4] ua[5] ua[6] ua[7] VGND
*.PININFO VPWR:I VGND:I ua[0]:B ena:I clk:I rst_n:I ua[1]:B ua[2]:B ua[3]:B ua[4]:B ua[5]:B ua[6]:B ua[7]:B uo_out[0]:O
*+ uo_out[1]:O uo_out[2]:O uo_out[3]:O uo_out[4]:O uo_out[5]:O uo_out[6]:O uo_out[7]:O ui_in[0]:I ui_in[1]:I ui_in[2]:I ui_in[3]:I ui_in[4]:I
*+ ui_in[5]:I ui_in[6]:I ui_in[7]:I uio_in[0]:I uio_in[1]:I uio_in[2]:I uio_in[3]:I uio_in[4]:I uio_in[5]:I uio_in[6]:I uio_in[7]:I
*+ uio_out[0]:O uio_out[1]:O uio_out[2]:O uio_out[3]:O uio_out[4]:O uio_out[5]:O uio_out[6]:O uio_out[7]:O uio_oe[0]:O uio_oe[1]:O uio_oe[2]:O
*+ uio_oe[3]:O uio_oe[4]:O uio_oe[5]:O uio_oe[6]:O uio_oe[7]:O
* noconn ua[2]
* noconn ua[3]
* noconn ua[4]
* noconn ua[5]
* noconn ua[6]
* noconn ua[7]
* noconn rst_n
* noconn clk
* noconn uio_in[0]
* noconn uio_in[1]
* noconn uio_in[2]
* noconn uio_in[3]
* noconn uio_in[4]
* noconn uio_in[5]
* noconn uio_in[6]
* noconn uio_in[7]
xdac VPWR dac_int ui_in[2] ui_in[1] ui_in[0] VGND dac
xringosc VPWR ro_int ui_in[6] VGND ringosc
* noconn ena
xtgro VPWR ua[0] ro_int ui_in[5] VGND tg
xtgdac VPWR ua[1] dac_int ui_in[3] VGND tg
xtgbyp VPWR ua[0] ua[1] ui_in[7] VGND tg
* noconn ui_in[4]
* noconn uo_out[7]
* noconn uo_out[6]
* noconn uo_out[5]
* noconn uo_out[4]
* noconn uo_out[3]
* noconn uo_out[2]
* noconn uo_out[1]
* noconn uo_out[0]
* noconn uio_out[7]
* noconn uio_out[6]
* noconn uio_out[5]
* noconn uio_out[4]
* noconn uio_out[3]
* noconn uio_out[2]
* noconn uio_out[1]
* noconn uio_out[0]
* noconn uio_oe[7]
* noconn uio_oe[0]
* noconn uio_oe[1]
* noconn uio_oe[2]
* noconn uio_oe[3]
* noconn uio_oe[4]
* noconn uio_oe[5]
* noconn uio_oe[6]
.ends

* expanding   symbol:  dac.sym # of pins=6
** sym_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/dac.sym
** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/dac.sch
.subckt dac vdd vout in2 in1 in0 vss
*.PININFO vdd:I vss:I vout:O in0:I in1:I in2:I
xdrv_b2 vdd in2 v2 vss dac_drv
xdrv_b1 vdd in1 v1 vss dac_drv
xdrv_b0 vdd in0 v0 vss dac_drv
XR1 net6 vout vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
xdrv_dummy vdd vss net4 vss dac_drv
XR2 net1 v2 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR3 vout net1 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
.save v(vout)
.save v(v2)
.save v(v1)
.save v(v0)
XR4 net5 net6 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR5 net7 v1 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR6 net6 net7 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR8 net2 v0 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR9 net5 net2 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR10 net3 net4 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR11 net5 net3 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XRdummy1 vss vss vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XRdummy2 vss vss vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
.ends


* expanding   symbol:  ringosc.sym # of pins=4
** sym_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc.sym
** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc.sch
.subckt ringosc vdd clk_out ena vss
*.PININFO vdd:I vss:I clk_out:O ena:I
.save v(ph1)
.save v(ph2)
.save v(ph3)
xro1 vdd ena ph1 ph2 vss ringosc_delay
xro2 vdd vdd ph2 ph3 vss ringosc_delay
xro3 vdd vdd ph3 ph1 vss ringosc_delay
xbuf1 vdd ph1 net1 vss ringosc_buf
xbuf2 vdd ph2 net2 vss ringosc_buf
xbuf3 vdd ph3 clk_out vss ringosc_buf
* noconn #net1
* noconn #net2
.save v(ena)
.ends


* expanding   symbol:  tg.sym # of pins=5
** sym_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/tg.sym
** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/tg.sch
.subckt tg vdd s1 s2 tgon vss
*.PININFO vdd:I vss:I tgon:I s2:B s1:B
XM3 s1 tgon s2 vss sky130_fd_pr__nfet_01v8 L=0.5 W=10 nf=1 m=1
XM4A s1 tgon_n s2 vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 m=1
XM4B s1 tgon_n s2 vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 m=1
XM1 tgon_n tgon vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM2 tgon_n tgon vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 m=1
.ends


* expanding   symbol:  dac_drv.sym # of pins=4
** sym_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/dac_drv.sym
** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/dac_drv.sch
.subckt dac_drv vdd in out vss
*.PININFO vdd:I vss:I in:I out:O
XM1 net1 in vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 m=1
XM2A net1 in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
XM4A out net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
XM3 out net1 vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 m=1
XM2B net1 in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
XM4B out net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
.ends


* expanding   symbol:  ringosc_delay.sym # of pins=5
** sym_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc_delay.sym
** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc_delay.sch
.subckt ringosc_delay vdd ena in out vss
*.PININFO vdd:I vss:I in:I out:O ena:I
XM1 out in vdd vdd sky130_fd_pr__pfet_01v8 L=10 W=0.5 nf=1 m=1
XM2A out in net1 vss sky130_fd_pr__nfet_01v8 L=10 W=0.5 nf=1 m=1
XMcap1 vss out vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=1 m=1
XMcap2 vdd out vdd vdd sky130_fd_pr__pfet_01v8 L=2 W=10 nf=1 m=1
XM2B net1 in vss vss sky130_fd_pr__nfet_01v8 L=10 W=0.5 nf=1 m=1
XMpowerdn in ena vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 m=1
.ends


* expanding   symbol:  ringosc_buf.sym # of pins=4
** sym_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc_buf.sym
** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc_buf.sch
.subckt ringosc_buf vdd in out vss
*.PININFO vdd:I vss:I in:I out:O
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=10 nf=1 m=1
XM2A out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 m=1
XM2B out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 m=1
.ends

.end
