** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/dac.sch
.subckt dac vdd vout in2 in1 in0 vss
*.PININFO vdd:I vss:I vout:O in0:I in1:I in2:I
xdrv_b2 vdd in2 v2 vss dac_drv
xdrv_b1 vdd in1 v1 vss dac_drv
xdrv_b0 vdd in0 v0 vss dac_drv
XR1 net6 vout vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
xdrv_dummy vdd vss net4 vss dac_drv
XR2 net1 v2 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR3 vout net1 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
.save v(vout)
.save v(v2)
.save v(v1)
.save v(v0)
XR4 net5 net6 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR5 net7 v1 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR6 net6 net7 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR8 net2 v0 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR9 net5 net2 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR10 net3 net4 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XR11 net5 net3 vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XRdummy1 vss vss vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
XRdummy2 vss vss vss sky130_fd_pr__res_xhigh_po_0p35 L=1.4 mult=1 m=1
.ends

* expanding   symbol:  dac_drv.sym # of pins=4
** sym_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/dac_drv.sym
** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/dac_drv.sch
.subckt dac_drv vdd in out vss
*.PININFO vdd:I vss:I in:I out:O
XM1 net1 in vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 m=1
XM2A net1 in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
XM4A out net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
XM3 out net1 vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 m=1
XM2B net1 in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
XM4B out net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
.ends

.end
