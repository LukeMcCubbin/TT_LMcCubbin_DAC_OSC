** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/dac_drv.sch
.subckt dac_drv vdd in out vss
*.PININFO vdd:I vss:I in:I out:O
XM1 net1 in vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 m=1
XM2A net1 in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
XM4A out net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
XM3 out net1 vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=1 m=1
XM2B net1 in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
XM4B out net1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=1 m=1
.ends
.end
