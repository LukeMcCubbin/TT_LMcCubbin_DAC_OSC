magic
tech sky130A
magscale 1 2
timestamp 1760644699
<< error_p >>
rect -1356 34 -1218 36
rect -1122 34 -984 36
rect -888 34 -750 36
rect -654 34 -516 36
rect -420 34 -282 36
rect -186 34 -48 36
rect 48 34 186 36
rect 282 34 420 36
rect 516 34 654 36
rect 750 34 888 36
rect 984 34 1122 36
rect 1218 34 1356 36
<< pwell >>
rect -1522 -632 1522 632
<< psubdiff >>
rect -1486 562 -1390 596
rect 1390 562 1486 596
rect -1486 500 -1452 562
rect 1452 500 1486 562
rect -1486 -562 -1452 -500
rect 1452 -562 1486 -500
rect -1486 -596 -1390 -562
rect 1390 -596 1486 -562
<< psubdiffcont >>
rect -1390 562 1390 596
rect -1486 -500 -1452 500
rect 1452 -500 1486 500
rect -1390 -596 1390 -562
<< xpolycontact >>
rect -1356 34 -1218 466
rect -1356 -466 -1218 -34
rect -1122 34 -984 466
rect -1122 -466 -984 -34
rect -888 34 -750 466
rect -888 -466 -750 -34
rect -654 34 -516 466
rect -654 -466 -516 -34
rect -420 34 -282 466
rect -420 -466 -282 -34
rect -186 34 -48 466
rect -186 -466 -48 -34
rect 48 34 186 466
rect 48 -466 186 -34
rect 282 34 420 466
rect 282 -466 420 -34
rect 516 34 654 466
rect 516 -466 654 -34
rect 750 34 888 466
rect 750 -466 888 -34
rect 984 34 1122 466
rect 984 -466 1122 -34
rect 1218 34 1356 466
rect 1218 -466 1356 -34
<< ppolyres >>
rect -1356 -34 -1218 34
rect -1122 -34 -984 34
rect -888 -34 -750 34
rect -654 -34 -516 34
rect -420 -34 -282 34
rect -186 -34 -48 34
rect 48 -34 186 34
rect 282 -34 420 34
rect 516 -34 654 34
rect 750 -34 888 34
rect 984 -34 1122 34
rect 1218 -34 1356 34
<< locali >>
rect -1486 562 -1390 596
rect 1390 562 1486 596
rect -1486 500 -1452 562
rect 1452 500 1486 562
rect -1486 -562 -1452 -500
rect 1452 -562 1486 -500
rect -1486 -596 -1390 -562
rect 1390 -596 1486 -562
<< viali >>
rect -1340 51 -1234 448
rect -1106 51 -1000 448
rect -872 51 -766 448
rect -638 51 -532 448
rect -404 51 -298 448
rect -170 51 -64 448
rect 64 51 170 448
rect 298 51 404 448
rect 532 51 638 448
rect 766 51 872 448
rect 1000 51 1106 448
rect 1234 51 1340 448
rect -1340 -448 -1234 -51
rect -1106 -448 -1000 -51
rect -872 -448 -766 -51
rect -638 -448 -532 -51
rect -404 -448 -298 -51
rect -170 -448 -64 -51
rect 64 -448 170 -51
rect 298 -448 404 -51
rect 532 -448 638 -51
rect 766 -448 872 -51
rect 1000 -448 1106 -51
rect 1234 -448 1340 -51
<< metal1 >>
rect -1346 448 -1228 460
rect -1346 51 -1340 448
rect -1234 51 -1228 448
rect -1346 39 -1228 51
rect -1112 448 -994 460
rect -1112 51 -1106 448
rect -1000 51 -994 448
rect -1112 39 -994 51
rect -878 448 -760 460
rect -878 51 -872 448
rect -766 51 -760 448
rect -878 39 -760 51
rect -644 448 -526 460
rect -644 51 -638 448
rect -532 51 -526 448
rect -644 39 -526 51
rect -410 448 -292 460
rect -410 51 -404 448
rect -298 51 -292 448
rect -410 39 -292 51
rect -176 448 -58 460
rect -176 51 -170 448
rect -64 51 -58 448
rect -176 39 -58 51
rect 58 448 176 460
rect 58 51 64 448
rect 170 51 176 448
rect 58 39 176 51
rect 292 448 410 460
rect 292 51 298 448
rect 404 51 410 448
rect 292 39 410 51
rect 526 448 644 460
rect 526 51 532 448
rect 638 51 644 448
rect 526 39 644 51
rect 760 448 878 460
rect 760 51 766 448
rect 872 51 878 448
rect 760 39 878 51
rect 994 448 1112 460
rect 994 51 1000 448
rect 1106 51 1112 448
rect 994 39 1112 51
rect 1228 448 1346 460
rect 1228 51 1234 448
rect 1340 51 1346 448
rect 1228 39 1346 51
rect -1346 -51 -1228 -39
rect -1346 -448 -1340 -51
rect -1234 -448 -1228 -51
rect -1346 -460 -1228 -448
rect -1112 -51 -994 -39
rect -1112 -448 -1106 -51
rect -1000 -448 -994 -51
rect -1112 -460 -994 -448
rect -878 -51 -760 -39
rect -878 -448 -872 -51
rect -766 -448 -760 -51
rect -878 -460 -760 -448
rect -644 -51 -526 -39
rect -644 -448 -638 -51
rect -532 -448 -526 -51
rect -644 -460 -526 -448
rect -410 -51 -292 -39
rect -410 -448 -404 -51
rect -298 -448 -292 -51
rect -410 -460 -292 -448
rect -176 -51 -58 -39
rect -176 -448 -170 -51
rect -64 -448 -58 -51
rect -176 -460 -58 -448
rect 58 -51 176 -39
rect 58 -448 64 -51
rect 170 -448 176 -51
rect 58 -460 176 -448
rect 292 -51 410 -39
rect 292 -448 298 -51
rect 404 -448 410 -51
rect 292 -460 410 -448
rect 526 -51 644 -39
rect 526 -448 532 -51
rect 638 -448 644 -51
rect 526 -460 644 -448
rect 760 -51 878 -39
rect 760 -448 766 -51
rect 872 -448 878 -51
rect 760 -460 878 -448
rect 994 -51 1112 -39
rect 994 -448 1000 -51
rect 1106 -448 1112 -51
rect 994 -460 1112 -448
rect 1228 -51 1346 -39
rect 1228 -448 1234 -51
rect 1340 -448 1346 -51
rect 1228 -460 1346 -448
<< properties >>
string FIXED_BBOX -1469 -579 1469 579
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 0.50 m 1 nx 12 wmin 0.690 lmin 0.50 rho 319.8 val 1.57k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
