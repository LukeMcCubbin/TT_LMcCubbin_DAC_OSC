magic
tech sky130A
magscale 1 2
timestamp 1759510403
<< pwell >>
rect -201 -722 201 722
<< psubdiff >>
rect -165 652 -69 686
rect 69 652 165 686
rect -165 590 -131 652
rect 131 590 165 652
rect -165 -652 -131 -590
rect 131 -652 165 -590
rect -165 -686 -69 -652
rect 69 -686 165 -652
<< psubdiffcont >>
rect -69 652 69 686
rect -165 -590 -131 590
rect 131 -590 165 590
rect -69 -686 69 -652
<< xpolycontact >>
rect -35 124 35 556
rect -35 -556 35 -124
<< xpolyres >>
rect -35 -124 35 124
<< locali >>
rect -165 652 -69 686
rect 69 652 165 686
rect -165 590 -131 652
rect 131 590 165 652
rect -165 -652 -131 -590
rect 131 -652 165 -590
rect -165 -686 -69 -652
rect 69 -686 165 -652
<< viali >>
rect -19 141 19 538
rect -19 -538 19 -141
<< metal1 >>
rect -25 538 25 550
rect -25 141 -19 538
rect 19 141 25 538
rect -25 129 25 141
rect -25 -141 25 -129
rect -25 -538 -19 -141
rect 19 -538 25 -141
rect -25 -550 25 -538
<< properties >>
string FIXED_BBOX -148 -669 148 669
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.4 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 9.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
