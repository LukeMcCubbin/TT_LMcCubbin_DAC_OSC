magic
tech sky130A
timestamp 1759510403
<< pwell >>
rect -598 -130 598 130
<< nmos >>
rect -500 -25 500 25
<< ndiff >>
rect -529 19 -500 25
rect -529 -19 -523 19
rect -506 -19 -500 19
rect -529 -25 -500 -19
rect 500 19 529 25
rect 500 -19 506 19
rect 523 -19 529 19
rect 500 -25 529 -19
<< ndiffc >>
rect -523 -19 -506 19
rect 506 -19 523 19
<< psubdiff >>
rect -580 95 -532 112
rect 532 95 580 112
rect -580 64 -563 95
rect 563 64 580 95
rect -580 -95 -563 -64
rect 563 -95 580 -64
rect -580 -112 -532 -95
rect 532 -112 580 -95
<< psubdiffcont >>
rect -532 95 532 112
rect -580 -64 -563 64
rect 563 -64 580 64
rect -532 -112 532 -95
<< poly >>
rect -500 61 500 69
rect -500 44 -492 61
rect 492 44 500 61
rect -500 25 500 44
rect -500 -44 500 -25
rect -500 -61 -492 -44
rect 492 -61 500 -44
rect -500 -69 500 -61
<< polycont >>
rect -492 44 492 61
rect -492 -61 492 -44
<< locali >>
rect -580 95 -532 112
rect 532 95 580 112
rect -580 64 -563 95
rect 563 64 580 95
rect -500 44 -492 61
rect 492 44 500 61
rect -523 19 -506 27
rect -523 -27 -506 -19
rect 506 19 523 27
rect 506 -27 523 -19
rect -500 -61 -492 -44
rect 492 -61 500 -44
rect -580 -95 -563 -64
rect 563 -95 580 -64
rect -580 -112 -532 -95
rect 532 -112 580 -95
<< viali >>
rect -492 44 492 61
rect -523 -19 -506 19
rect 506 -19 523 19
rect -492 -61 492 -44
<< metal1 >>
rect -498 61 498 64
rect -498 44 -492 61
rect 492 44 498 61
rect -498 41 498 44
rect -526 19 -503 25
rect -526 -19 -523 19
rect -506 -19 -503 19
rect -526 -25 -503 -19
rect 503 19 526 25
rect 503 -19 506 19
rect 523 -19 526 19
rect 503 -25 526 -19
rect -498 -44 498 -41
rect -498 -61 -492 -44
rect 492 -61 498 -44
rect -498 -64 498 -61
<< properties >>
string FIXED_BBOX -571 -103 571 103
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 10.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
