magic
tech sky130A
magscale 1 2
timestamp 1760719168
<< pwell >>
rect -4487 -250 -1443 1052
<< psubdiff >>
rect -4451 982 -4355 1016
rect -1575 982 -1479 1016
rect -4451 920 -4417 982
rect -1513 920 -1479 982
rect -4451 -180 -4417 -118
rect -1513 -180 -1479 -118
rect -4451 -214 -4355 -180
rect -1575 -214 -1479 -180
<< psubdiffcont >>
rect -4355 982 -1575 1016
rect -4451 -118 -4417 920
rect -1513 -118 -1479 920
rect -4355 -214 -1575 -180
<< xpolycontact >>
rect -4321 454 -4183 886
rect -4321 -84 -4183 348
rect -4087 454 -3949 886
rect -4087 -84 -3949 348
rect -3853 454 -3715 886
rect -3853 -84 -3715 348
rect -3619 454 -3481 886
rect -3619 -84 -3481 348
rect -3385 454 -3247 886
rect -3385 -84 -3247 348
rect -3151 454 -3013 886
rect -3151 -84 -3013 348
rect -2917 454 -2779 886
rect -2917 -84 -2779 348
rect -2683 454 -2545 886
rect -2683 -84 -2545 348
rect -2449 454 -2311 886
rect -2449 -84 -2311 348
rect -2215 454 -2077 886
rect -2215 -84 -2077 348
rect -1981 454 -1843 886
rect -1981 -84 -1843 348
rect -1747 454 -1609 886
rect -1747 -84 -1609 348
<< ppolyres >>
rect -4321 348 -4183 454
rect -4087 348 -3949 454
rect -3853 348 -3715 454
rect -3619 348 -3481 454
rect -3385 348 -3247 454
rect -3151 348 -3013 454
rect -2917 348 -2779 454
rect -2683 348 -2545 454
rect -2449 348 -2311 454
rect -2215 348 -2077 454
rect -1981 348 -1843 454
rect -1747 348 -1609 454
<< locali >>
rect -4451 982 -4355 1016
rect -1575 982 -1479 1016
rect -4451 920 -4417 982
rect -1513 920 -1479 982
rect -4451 -180 -4417 -118
rect -1513 -180 -1479 -118
rect -4451 -214 -4355 -180
rect -1575 -214 -1479 -180
<< properties >>
string FIXED_BBOX -1469 -598 1469 598
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 0.69 m 1 nx 12 wmin 0.690 lmin 0.50 rho 319.8 val 884.495 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
