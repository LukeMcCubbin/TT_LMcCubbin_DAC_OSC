magic
tech sky130A
magscale 1 2
timestamp 1760463315
<< metal3 >>
rect 200 18111 9248 18112
rect 195 17713 201 18111
rect 599 17713 9248 18111
rect 200 17712 9248 17713
rect 9648 17712 9654 18112
rect 8409 1152 8807 1157
rect 8408 1151 17934 1152
rect 8408 753 8409 1151
rect 8807 753 17934 1151
rect 8408 752 17934 753
rect 18334 752 18340 1152
rect 8409 747 8807 752
<< via3 >>
rect 201 17713 599 18111
rect 9248 17712 9648 18112
rect 8409 753 8807 1151
rect 17934 752 18334 1152
<< metal4 >>
rect 200 18111 600 44152
rect 800 44082 1200 44152
rect 800 43422 1194 44082
rect 800 24716 1200 43422
rect 6134 41940 6194 45152
rect 4294 41880 6210 41940
rect 796 24316 2844 24716
rect 200 17713 201 18111
rect 599 17713 600 18111
rect 200 1000 600 17713
rect 800 1000 1200 24316
rect 2444 19204 2844 24316
rect 4294 22220 4354 41880
rect 6134 41862 6194 41880
rect 6686 41544 6746 45152
rect 4846 41484 6780 41544
rect 4846 22224 4906 41484
rect 6686 41462 6746 41484
rect 5398 41380 5458 41392
rect 7238 41380 7298 45152
rect 5398 41320 7298 41380
rect 5398 22220 5458 41320
rect 7238 41316 7298 41320
rect 5950 41190 6010 41198
rect 7790 41190 7850 45152
rect 5950 41130 7850 41190
rect 5950 22238 6010 41130
rect 6502 41010 6562 41028
rect 8342 41010 8402 45152
rect 6502 40950 8404 41010
rect 6502 22224 6562 40950
rect 8342 40918 8402 40950
rect 8894 40846 8954 45152
rect 7054 40786 8956 40846
rect 7054 22224 7114 40786
rect 8894 40754 8954 40786
rect 9446 40608 9506 45152
rect 7606 40548 9510 40608
rect 7606 22208 7666 40548
rect 9446 40484 9506 40548
rect 9998 40188 10058 45152
rect 8156 40128 10058 40188
rect 8156 24340 8216 40128
rect 9998 40110 10058 40128
rect 8710 40028 8770 40036
rect 10550 40028 10610 45152
rect 8710 39968 10612 40028
rect 8156 24214 8218 24340
rect 8158 22224 8218 24214
rect 8710 22216 8770 39968
rect 10550 39928 10610 39968
rect 9262 39714 9322 39730
rect 11102 39714 11162 45152
rect 9262 39654 11162 39714
rect 9262 22216 9322 39654
rect 11102 39618 11162 39654
rect 9814 39334 9874 39350
rect 11654 39334 11714 45152
rect 9814 39274 11714 39334
rect 9814 22202 9874 39274
rect 11654 39218 11714 39274
rect 10366 38970 10426 38994
rect 12206 38970 12266 45152
rect 10366 38910 12266 38970
rect 10366 22212 10426 38910
rect 12206 38898 12266 38910
rect 12758 38582 12818 45152
rect 10918 38522 12820 38582
rect 10918 22226 10978 38522
rect 12758 38504 12818 38522
rect 13310 38322 13370 45152
rect 11470 38262 13370 38322
rect 11470 22218 11530 38262
rect 13310 38226 13370 38262
rect 13862 38020 13922 45152
rect 12022 37960 13924 38020
rect 12022 22208 12082 37960
rect 13862 37936 13922 37960
rect 14414 37694 14474 45152
rect 12574 37634 14474 37694
rect 12574 22200 12634 37634
rect 14966 37326 15026 45152
rect 13126 37266 15028 37326
rect 13126 22200 13186 37266
rect 14966 37260 15026 37266
rect 13678 36956 13738 36960
rect 15518 36956 15578 45152
rect 13678 36896 15580 36956
rect 13678 22164 13738 36896
rect 15518 36854 15578 36896
rect 16070 36526 16130 45152
rect 14230 36466 16132 36526
rect 14230 22208 14290 36466
rect 16070 36436 16130 36466
rect 16622 36158 16682 45152
rect 14782 36098 16684 36158
rect 14782 22184 14842 36098
rect 16622 36058 16682 36098
rect 17174 35856 17234 45152
rect 15334 35796 17234 35856
rect 15334 22218 15394 35796
rect 17174 35748 17234 35796
rect 17726 35358 17786 45152
rect 15902 35298 17788 35358
rect 15902 22190 15962 35298
rect 17726 35242 17786 35298
rect 16438 34772 16498 34818
rect 18278 34772 18338 45152
rect 16438 34712 18338 34772
rect 16438 22218 16498 34712
rect 18278 34706 18338 34712
rect 16990 34370 17050 34406
rect 18830 34370 18890 45152
rect 19382 44870 19442 45152
rect 19934 44870 19994 45152
rect 20486 44870 20546 45152
rect 21038 44870 21098 45152
rect 21590 44870 21650 45152
rect 22142 44870 22202 45152
rect 22694 44870 22754 45152
rect 23246 44870 23306 45152
rect 23798 36280 23858 45152
rect 16990 34310 18890 34370
rect 21958 36220 23858 36280
rect 16990 22148 17050 34310
rect 17542 22184 17602 22442
rect 21958 22172 22018 36220
rect 23798 36212 23858 36220
rect 24350 35826 24410 45152
rect 22510 35766 24438 35826
rect 22510 22172 22570 35766
rect 24902 35442 24962 45152
rect 25454 44896 25514 45152
rect 23062 35382 25002 35442
rect 23062 22200 23122 35382
rect 24902 35372 24962 35382
rect 26006 34714 26066 45152
rect 24166 34654 26080 34714
rect 24166 22154 24226 34654
rect 26006 34632 26066 34654
rect 26558 34276 26618 45152
rect 24718 34216 26628 34276
rect 24718 22146 24778 34216
rect 26558 34204 26618 34216
rect 27110 33820 27170 45152
rect 25270 33760 27176 33820
rect 25270 22182 25330 33760
rect 27110 33742 27170 33760
rect 27662 33364 27722 45152
rect 25822 33304 27732 33364
rect 25822 22182 25882 33304
rect 27662 33286 27722 33304
rect 28214 33016 28274 45152
rect 26374 32956 28276 33016
rect 26374 22224 26434 32956
rect 28214 32928 28274 32956
rect 28766 32646 28826 45152
rect 26926 32586 28826 32646
rect 26926 22210 26986 32586
rect 28766 32546 28826 32586
rect 29318 32264 29378 45152
rect 27478 32204 29378 32264
rect 27478 22204 27538 32204
rect 29318 32180 29378 32204
rect 2444 18804 8008 19204
rect 7608 1152 8008 18804
rect 9247 18112 9649 18113
rect 11132 18112 11548 18134
rect 9247 17712 9248 18112
rect 9648 17712 12964 18112
rect 9247 17711 9649 17712
rect 11132 17242 11548 17712
rect 11132 16508 12464 17242
rect 11148 16486 12464 16508
rect 17933 1152 18335 1153
rect 7608 1151 8808 1152
rect 7608 753 8409 1151
rect 8807 753 8808 1151
rect 7608 752 8808 753
rect 17933 752 17934 1152
rect 18334 752 20256 1152
rect 17933 751 18335 752
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 194 26678 200
rect 26160 14 26678 194
rect 26498 0 26678 14
rect 30362 0 30542 510
use tt_um_tt05_analog_test_cell  tt_um_tt05_analog_test_cell_0
timestamp 1760454724
transform 1 0 0 0 1 0
box 768 0 30594 22304
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel space 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
rlabel metal4 800 1000 1200 43422 1 VGND
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
