magic
tech sky130A
magscale 1 2
timestamp 1759510403
<< nwell >>
rect -1196 -269 1196 269
<< pmos >>
rect -1000 -50 1000 50
<< pdiff >>
rect -1058 38 -1000 50
rect -1058 -38 -1046 38
rect -1012 -38 -1000 38
rect -1058 -50 -1000 -38
rect 1000 38 1058 50
rect 1000 -38 1012 38
rect 1046 -38 1058 38
rect 1000 -50 1058 -38
<< pdiffc >>
rect -1046 -38 -1012 38
rect 1012 -38 1046 38
<< nsubdiff >>
rect -1160 199 -1064 233
rect 1064 199 1160 233
rect -1160 137 -1126 199
rect 1126 137 1160 199
rect -1160 -199 -1126 -137
rect 1126 -199 1160 -137
rect -1160 -233 -1064 -199
rect 1064 -233 1160 -199
<< nsubdiffcont >>
rect -1064 199 1064 233
rect -1160 -137 -1126 137
rect 1126 -137 1160 137
rect -1064 -233 1064 -199
<< poly >>
rect -1000 131 1000 147
rect -1000 97 -984 131
rect 984 97 1000 131
rect -1000 50 1000 97
rect -1000 -97 1000 -50
rect -1000 -131 -984 -97
rect 984 -131 1000 -97
rect -1000 -147 1000 -131
<< polycont >>
rect -984 97 984 131
rect -984 -131 984 -97
<< locali >>
rect -1160 199 -1064 233
rect 1064 199 1160 233
rect -1160 137 -1126 199
rect 1126 137 1160 199
rect -1000 97 -984 131
rect 984 97 1000 131
rect -1046 38 -1012 54
rect -1046 -54 -1012 -38
rect 1012 38 1046 54
rect 1012 -54 1046 -38
rect -1000 -131 -984 -97
rect 984 -131 1000 -97
rect -1160 -199 -1126 -137
rect 1126 -199 1160 -137
rect -1160 -233 -1064 -199
rect 1064 -233 1160 -199
<< viali >>
rect -984 97 984 131
rect -1046 -38 -1012 38
rect 1012 -38 1046 38
rect -984 -131 984 -97
<< metal1 >>
rect -996 131 996 137
rect -996 97 -984 131
rect 984 97 996 131
rect -996 91 996 97
rect -1052 38 -1006 50
rect -1052 -38 -1046 38
rect -1012 -38 -1006 38
rect -1052 -50 -1006 -38
rect 1006 38 1052 50
rect 1006 -38 1012 38
rect 1046 -38 1052 38
rect 1006 -50 1052 -38
rect -996 -97 996 -91
rect -996 -131 -984 -97
rect 984 -131 996 -97
rect -996 -137 996 -131
<< properties >>
string FIXED_BBOX -1143 -216 1143 216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 10.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
