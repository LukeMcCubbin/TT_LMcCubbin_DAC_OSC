** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc.sch
.subckt ringosc vdd clk_out ena vss
*.PININFO vdd:I vss:I clk_out:O ena:I
.save v(ph1)
.save v(ph2)
.save v(ph3)
xro1 vdd ena ph1 ph2 vss ringosc_delay
xro2 vdd vdd ph2 ph3 vss ringosc_delay
xro3 vdd vdd ph3 ph1 vss ringosc_delay
xbuf1 vdd ph1 net1 vss ringosc_buf
xbuf2 vdd ph2 net2 vss ringosc_buf
xbuf3 vdd ph3 clk_out vss ringosc_buf
* noconn #net1
* noconn #net2
.save v(ena)
.ends

* expanding   symbol:  ringosc_delay.sym # of pins=5
** sym_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc_delay.sym
** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc_delay.sch
.subckt ringosc_delay vdd ena in out vss
*.PININFO vdd:I vss:I in:I out:O ena:I
XM1 out in vdd vdd sky130_fd_pr__pfet_01v8 L=10 W=0.5 nf=1 m=1
XM2A out in net1 vss sky130_fd_pr__nfet_01v8 L=10 W=0.5 nf=1 m=1
XMcap1 vss out vss vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=1 m=1
XMcap2 vdd out vdd vdd sky130_fd_pr__pfet_01v8 L=2 W=10 nf=1 m=1
XM2B net1 in vss vss sky130_fd_pr__nfet_01v8 L=10 W=0.5 nf=1 m=1
XMpowerdn in ena vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 m=1
.ends


* expanding   symbol:  ringosc_buf.sym # of pins=4
** sym_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc_buf.sym
** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/ringosc_buf.sch
.subckt ringosc_buf vdd in out vss
*.PININFO vdd:I vss:I in:I out:O
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=10 nf=1 m=1
XM2A out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 m=1
XM2B out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 m=1
.ends

.end
