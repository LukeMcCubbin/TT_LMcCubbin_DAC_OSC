magic
tech sky130A
timestamp 1759510403
<< pwell >>
rect -198 -605 198 605
<< nmos >>
rect -100 -500 100 500
<< ndiff >>
rect -129 494 -100 500
rect -129 -494 -123 494
rect -106 -494 -100 494
rect -129 -500 -100 -494
rect 100 494 129 500
rect 100 -494 106 494
rect 123 -494 129 494
rect 100 -500 129 -494
<< ndiffc >>
rect -123 -494 -106 494
rect 106 -494 123 494
<< psubdiff >>
rect -180 570 -132 587
rect 132 570 180 587
rect -180 539 -163 570
rect 163 539 180 570
rect -180 -570 -163 -539
rect 163 -570 180 -539
rect -180 -587 -132 -570
rect 132 -587 180 -570
<< psubdiffcont >>
rect -132 570 132 587
rect -180 -539 -163 539
rect 163 -539 180 539
rect -132 -587 132 -570
<< poly >>
rect -100 536 100 544
rect -100 519 -92 536
rect 92 519 100 536
rect -100 500 100 519
rect -100 -519 100 -500
rect -100 -536 -92 -519
rect 92 -536 100 -519
rect -100 -544 100 -536
<< polycont >>
rect -92 519 92 536
rect -92 -536 92 -519
<< locali >>
rect -180 570 -132 587
rect 132 570 180 587
rect -180 539 -163 570
rect 163 539 180 570
rect -100 519 -92 536
rect 92 519 100 536
rect -123 494 -106 502
rect -123 -502 -106 -494
rect 106 494 123 502
rect 106 -502 123 -494
rect -100 -536 -92 -519
rect 92 -536 100 -519
rect -180 -570 -163 -539
rect 163 -570 180 -539
rect -180 -587 -132 -570
rect 132 -587 180 -570
<< viali >>
rect -92 519 92 536
rect -123 -494 -106 494
rect 106 -494 123 494
rect -92 -536 92 -519
<< metal1 >>
rect -98 536 98 539
rect -98 519 -92 536
rect 92 519 98 536
rect -98 516 98 519
rect -126 494 -103 500
rect -126 -494 -123 494
rect -106 -494 -103 494
rect -126 -500 -103 -494
rect 103 494 126 500
rect 103 -494 106 494
rect 123 -494 126 494
rect 103 -500 126 -494
rect -98 -519 98 -516
rect -98 -536 -92 -519
rect 92 -536 98 -519
rect -98 -539 98 -536
<< properties >>
string FIXED_BBOX -171 -578 171 578
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
