magic
tech sky130A
magscale 1 2
timestamp 1760727663
use res_str  sky130_fd_pr__res_high_po_0p69_AWHN5X_0
timestamp 1760719168
transform 1 0 355 0 1 -140
box -4487 -250 -1443 1052
<< properties >>
string FIXED_BBOX -1060 -684 1060 684
<< end >>
