magic
tech sky130A
magscale 1 2
timestamp 1761151864
<< pwell >>
rect -1522 -651 1522 651
<< psubdiff >>
rect -1486 581 -1390 615
rect 1390 581 1486 615
rect -1486 -581 -1452 581
rect 1452 -581 1486 581
rect -1486 -615 -1390 -581
rect 1390 -615 1486 -581
<< psubdiffcont >>
rect -1390 581 1390 615
rect -1390 -615 1390 -581
<< xpolycontact >>
rect -1356 53 -1218 485
rect -1356 -485 -1218 -53
rect -1122 53 -984 485
rect -1122 -485 -984 -53
rect -888 53 -750 485
rect -888 -485 -750 -53
rect -654 53 -516 485
rect -654 -485 -516 -53
rect -420 53 -282 485
rect -420 -485 -282 -53
rect -186 53 -48 485
rect -186 -485 -48 -53
rect 48 53 186 485
rect 48 -485 186 -53
rect 282 53 420 485
rect 282 -485 420 -53
rect 516 53 654 485
rect 516 -485 654 -53
rect 750 53 888 485
rect 750 -485 888 -53
rect 984 53 1122 485
rect 984 -485 1122 -53
rect 1218 53 1356 485
rect 1218 -485 1356 -53
<< ppolyres >>
rect -1356 -53 -1218 53
rect -1122 -53 -984 53
rect -888 -53 -750 53
rect -654 -53 -516 53
rect -420 -53 -282 53
rect -186 -53 -48 53
rect 48 -53 186 53
rect 282 -53 420 53
rect 516 -53 654 53
rect 750 -53 888 53
rect 984 -53 1122 53
rect 1218 -53 1356 53
<< locali >>
rect -1406 581 -1390 615
rect 1390 581 1406 615
rect -1406 -615 -1390 -581
rect 1390 -615 1406 -581
<< viali >>
rect -1340 70 -1234 467
rect -1106 70 -1000 467
rect -872 70 -766 467
rect -638 70 -532 467
rect -404 70 -298 467
rect -170 70 -64 467
rect 64 70 170 467
rect 298 70 404 467
rect 532 70 638 467
rect 766 70 872 467
rect 1000 70 1106 467
rect 1234 70 1340 467
rect -1340 -467 -1234 -70
rect -1106 -467 -1000 -70
rect -872 -467 -766 -70
rect -638 -467 -532 -70
rect -404 -467 -298 -70
rect -170 -467 -64 -70
rect 64 -467 170 -70
rect 298 -467 404 -70
rect 532 -467 638 -70
rect 766 -467 872 -70
rect 1000 -467 1106 -70
rect 1234 -467 1340 -70
<< metal1 >>
rect -1346 467 -1228 479
rect -1346 70 -1340 467
rect -1234 70 -1228 467
rect -1346 58 -1228 70
rect -1112 467 -994 479
rect -1112 70 -1106 467
rect -1000 70 -994 467
rect -1112 58 -994 70
rect -878 467 -760 479
rect -878 70 -872 467
rect -766 70 -760 467
rect -878 58 -760 70
rect -644 467 -526 479
rect -644 70 -638 467
rect -532 70 -526 467
rect -644 58 -526 70
rect -410 467 -292 479
rect -410 70 -404 467
rect -298 70 -292 467
rect -410 58 -292 70
rect -176 467 -58 479
rect -176 70 -170 467
rect -64 70 -58 467
rect -176 58 -58 70
rect 58 467 176 479
rect 58 70 64 467
rect 170 70 176 467
rect 58 58 176 70
rect 292 467 410 479
rect 292 70 298 467
rect 404 70 410 467
rect 292 58 410 70
rect 526 467 644 479
rect 526 70 532 467
rect 638 70 644 467
rect 526 58 644 70
rect 760 467 878 479
rect 760 70 766 467
rect 872 70 878 467
rect 760 58 878 70
rect 994 467 1112 479
rect 994 70 1000 467
rect 1106 70 1112 467
rect 994 58 1112 70
rect 1228 467 1346 479
rect 1228 70 1234 467
rect 1340 70 1346 467
rect 1228 58 1346 70
rect -1346 -70 -1228 -58
rect -1346 -467 -1340 -70
rect -1234 -467 -1228 -70
rect -1346 -479 -1228 -467
rect -1112 -70 -994 -58
rect -1112 -467 -1106 -70
rect -1000 -467 -994 -70
rect -1112 -479 -994 -467
rect -878 -70 -760 -58
rect -878 -467 -872 -70
rect -766 -467 -760 -70
rect -878 -479 -760 -467
rect -644 -70 -526 -58
rect -644 -467 -638 -70
rect -532 -467 -526 -70
rect -644 -479 -526 -467
rect -410 -70 -292 -58
rect -410 -467 -404 -70
rect -298 -467 -292 -70
rect -410 -479 -292 -467
rect -176 -70 -58 -58
rect -176 -467 -170 -70
rect -64 -467 -58 -70
rect -176 -479 -58 -467
rect 58 -70 176 -58
rect 58 -467 64 -70
rect 170 -467 176 -70
rect 58 -479 176 -467
rect 292 -70 410 -58
rect 292 -467 298 -70
rect 404 -467 410 -70
rect 292 -479 410 -467
rect 526 -70 644 -58
rect 526 -467 532 -70
rect 638 -467 644 -70
rect 526 -479 644 -467
rect 760 -70 878 -58
rect 760 -467 766 -70
rect 872 -467 878 -70
rect 760 -479 878 -467
rect 994 -70 1112 -58
rect 994 -467 1000 -70
rect 1106 -467 1112 -70
rect 994 -479 1112 -467
rect 1228 -70 1346 -58
rect 1228 -467 1234 -70
rect 1340 -467 1346 -70
rect 1228 -479 1346 -467
<< properties >>
string FIXED_BBOX -1469 -598 1469 598
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 0.690 m 1 nx 12 wmin 0.690 lmin 0.50 rho 319.8 val 884.495 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 0 grc 0 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 0 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
