magic
tech sky130A
timestamp 1760644699
<< error_p >>
rect -678 17 -609 18
rect -561 17 -492 18
rect -444 17 -375 18
rect -327 17 -258 18
rect -210 17 -141 18
rect -93 17 -24 18
rect 24 17 93 18
rect 141 17 210 18
rect 258 17 327 18
rect 375 17 444 18
rect 492 17 561 18
rect 609 17 678 18
<< pwell >>
rect -761 -316 761 316
<< psubdiff >>
rect -743 281 -695 298
rect 695 281 743 298
rect -743 250 -726 281
rect 726 250 743 281
rect -743 -281 -726 -250
rect 726 -281 743 -250
rect -743 -298 -695 -281
rect 695 -298 743 -281
<< psubdiffcont >>
rect -695 281 695 298
rect -743 -250 -726 250
rect 726 -250 743 250
rect -695 -298 695 -281
<< xpolycontact >>
rect -678 17 -609 233
rect -678 -233 -609 -17
rect -561 17 -492 233
rect -561 -233 -492 -17
rect -444 17 -375 233
rect -444 -233 -375 -17
rect -327 17 -258 233
rect -327 -233 -258 -17
rect -210 17 -141 233
rect -210 -233 -141 -17
rect -93 17 -24 233
rect -93 -233 -24 -17
rect 24 17 93 233
rect 24 -233 93 -17
rect 141 17 210 233
rect 141 -233 210 -17
rect 258 17 327 233
rect 258 -233 327 -17
rect 375 17 444 233
rect 375 -233 444 -17
rect 492 17 561 233
rect 492 -233 561 -17
rect 609 17 678 233
rect 609 -233 678 -17
<< ppolyres >>
rect -678 -17 -609 17
rect -561 -17 -492 17
rect -444 -17 -375 17
rect -327 -17 -258 17
rect -210 -17 -141 17
rect -93 -17 -24 17
rect 24 -17 93 17
rect 141 -17 210 17
rect 258 -17 327 17
rect 375 -17 444 17
rect 492 -17 561 17
rect 609 -17 678 17
<< locali >>
rect -743 281 -695 298
rect 695 281 743 298
rect -743 250 -726 281
rect 726 250 743 281
rect -743 -281 -726 -250
rect 726 -281 743 -250
rect -743 -298 -695 -281
rect 695 -298 743 -281
<< properties >>
string FIXED_BBOX -734 -289 734 289
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 0.50 m 1 nx 12 wmin 0.690 lmin 0.50 rho 319.8 val 796.434 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
