** sch_path: /home/ttuser/TT_LMcCubbin_DAC_OSC/xschem/tg.sch
.subckt tg vdd s1 s2 tgon vss
*.PININFO vdd:I vss:I tgon:I s2:B s1:B
XM3 s1 tgon s2 vss sky130_fd_pr__nfet_01v8 L=0.5 W=10 nf=1 m=1
XM4A s1 tgon_n s2 vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 m=1
XM4B s1 tgon_n s2 vdd sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=1 m=1
XM1 tgon_n tgon vss vss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM2 tgon_n tgon vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 m=1
.ends
.end
